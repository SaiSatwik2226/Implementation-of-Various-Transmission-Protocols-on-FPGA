//////////////////////////////////////////////////////////////////////
// File Downloaded from http://www.nandland.com
//////////////////////////////////////////////////////////////////////

// This testbench will exercise the UART RX.
// It sends out byte 0x37, and ensures the RX receives it correctly.
`timescale 1ns/10ps

module UART_RX_TB();

  // Testbench uses a 25 MHz clock (same as Go Board)
  // Want to interface to 115200 baud UART
  // 25000000 / 115200 = 217 Clocks Per Bit.
  parameter c_CLOCK_PERIOD_NS = 10;
  parameter c_CLKS_PER_BIT    = 868;
  parameter c_BIT_PERIOD      = 8680;
  
  reg Clock = 0;
  reg RX_Serial = 1;
  wire [7:0] w_RX_Byte;
  wire RX_Done;
  
  // Takes in input byte and serializes it 
  task UART_WRITE_BYTE;
    input [7:0] i_Data;
    integer     ii;
    begin
      
      // Send Start Bit
      RX_Serial <= 1'b0;
      #(c_BIT_PERIOD);
      //#1000;
      
		
      // Send Data Byte
      for (ii=0; ii<8; ii=ii+1)
        begin
          RX_Serial <= i_Data[ii];
          #(c_BIT_PERIOD);
        end
      
      // Send Stop Bit
      RX_Serial <= 1'b1;
      #(c_BIT_PERIOD);
     end
  endtask // UART_WRITE_BYTE
  
  
  UART_RX #(.CLKS_PER_BIT(c_CLKS_PER_BIT)) UART_RX_INST
     (.Clock(Clock),
	  .RX_Serial(RX_Serial),
     //.RX_Done_Out(RX_Done_Out),
	  .RX_Done(RX_Done),
     .RX_Bytes(w_RX_Byte));
  
  always
    #(c_CLOCK_PERIOD_NS/2) Clock <= !Clock;

  
  // Main Testing:
  initial
    begin
      // Send a command to the UART (exercise Rx)
      //@(posedge Clock);
      UART_WRITE_BYTE(8'h37);
      //@(posedge Clock);
            
      // Check that the correct command was received
      if (w_RX_Byte == 8'h37)
        $display("Test Passed - Correct Byte Received");
      else
        $display("Test Failed - Incorrect Byte Received");
    $finish();
    end
endmodule

